LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY output IS 
	port(
		hour_upper_in:IN STD_LOGIC_VECTOR(3 downto 0);
		hour_lower_in:IN STD_LOGIC_VECTOR(3 downto 0);
		min_upper_in:IN STD_LOGIC_VECTOR(3 downto 0);
		min_lower_in:IN STD_LOGIC_VECTOR(3 downto 0);
		sec_upper_in:IN STD_LOGIC_VECTOR(3 downto 0);
		sec_lower_in:IN STD_LOGIC_VECTOR(3 downto 0);
		
		switch:in STD_LOGIC_VECTOR(1 DOWNTO 0);
		state:IN STD_LOGIC;
		ctr:in STD_LOGIC_VECTOR(1 DOWNTO 0);
		clk:in std_logic;
		
		sec_lower_7_out:OUT STD_LOGIC_VECTOR(6 downto 0);
		hour_lower_out:OUT STD_LOGIC_VECTOR(3 downto 0);
		min_upper_out:OUT STD_LOGIC_VECTOR(3 downto 0);
		min_lower_out:OUT STD_LOGIC_VECTOR(3 downto 0);
		sec_upper_out:OUT STD_LOGIC_VECTOR(3 downto 0);
		hour_upper_out:OUT STD_LOGIC_VECTOR(3 downto 0)
		);
END output;

ARCHITECTURE arch OF output IS
	SIGNAL var : STD_LOGIC_VECTOR(6 downto 0);
	BEGIN
	PROCESS(sec_lower_in)
	BEGIN
		CASE sec_lower_in IS
		WHEN "0000" => 
			var <= "1111110";
		WHEN "0001" => 
			var <= "0110000";
		WHEN "0010" => 
			var <= "1101101";
		WHEN "0011" => 
			var <= "1111001";
		WHEN "0100" => 
			var <= "0110011";
		WHEN "0101" =>
			var <= "1011011";
		WHEN "0110" => 
			var <= "1011111";
		WHEN "0111" =>
			var <= "1110000";
		WHEN "1000" => 
			var <= "1111111";
		WHEN "1001" =>
			var <= "1111011";
		WHEN OTHERS =>
			var <= "0001000";
		END CASE;
	END PROCESS;
	

	sec_lower_7_out<=var;
	sec_upper_out<=sec_upper_in;
	
	--hour_lower_out<=hour_lower_in;
	--hour_upper_out<=hour_upper_in;
	--min_lower_out<=min_lower_in;		
	--min_upper_out<=min_upper_in;	
	
	process(state,switch,ctr)
	begin
		if(state='0')then	
            min_upper_out<=min_upper_in;
            min_lower_out<=min_lower_in;
			hour_lower_out<=hour_lower_in;
			hour_upper_out<=hour_upper_in;
		elsif(state='1')then
			case(switch)is
				when"00"=>
					hour_lower_out<=hour_lower_in;
					hour_upper_out<=hour_upper_in;
					min_lower_out<=min_lower_in;		
					min_upper_out<=min_upper_in;
				when"01"=>
					hour_lower_out<=hour_lower_in;
					hour_upper_out<=hour_upper_in;
					case(clk)is
						when '1'=>
						min_lower_out<="ZZZZ";		
						min_upper_out<="ZZZZ";
						when others=>
						min_lower_out<=min_lower_in;		
						min_upper_out<=min_upper_in;
					end case;
				when"10"=>
					min_lower_out<=min_lower_in;		
					min_upper_out<=min_upper_in;				
					case(clk)is
						when '1'=>
						hour_lower_out<="ZZZZ";
						hour_upper_out<="ZZZZ";
						when others=>
						hour_lower_out<=hour_lower_in;
						hour_upper_out<=hour_upper_in;
					end case;
				when others=>
									
					case(clk)is
						when '1'=>
						hour_lower_out<="ZZZZ";
						hour_upper_out<="ZZZZ";
						min_lower_out<="ZZZZ";		
						min_upper_out<="ZZZZ";
						when others=>
						min_lower_out<=min_lower_in;		
						min_upper_out<=min_upper_in;
						hour_lower_out<=hour_lower_in;
						hour_upper_out<=hour_upper_in;
					end case;
				end case;
			end if;
		end process;		
END arch;